module Restador(
	input logic a, 
	input logic b, 
	input logic cin, 
	output logic d, 
	output logic bo
);


endmodule
