library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FourBitAdder_FPGA is
    Port ( 
	 
			SW : in  STD_LOGIC_VECTOR (7 downto 0); 
			Cin : in  STD_LOGIC; 
			HEX : out STD_LOGIC_VECTOR (6 downto 0);
			Cout : out STD_LOGIC); 
			
	end FourBitAdder_FPGA;

architecture Behavioral of FourBitAdder_FPGA is
    component FourBitAdder
        Port ( 
				A : in  STD_LOGIC_VECTOR (3 downto 0);
				B : in  STD_LOGIC_VECTOR (3 downto 0);
				Cin : in  STD_LOGIC;
				Sum : out STD_LOGIC_VECTOR (3 downto 0);
				Cout : out STD_LOGIC);
				
    end component;

    signal A, B, Sum : STD_LOGIC_VECTOR (3 downto 0);
    
begin
    A <= SW(7 downto 4);
    B <= SW(3 downto 0);

    SUMADOR: FourBitAdder port map(A, B, Cin, Sum, Cout);

    -- Conversión del resultado a 7 segmentos
    process(Sum)
    begin
        case Sum is
		  
            when "0000" => HEX <= "1000000"; -- 0
            when "0001" => HEX <= "1111001"; -- 1
            when "0010" => HEX <= "0100100"; -- 2
            when "0011" => HEX <= "0110000"; -- 3
            when "0100" => HEX <= "0011001"; -- 4
            when "0101" => HEX <= "0010010"; -- 5
            when "0110" => HEX <= "0000010"; -- 6
            when "0111" => HEX <= "1111000"; -- 7
            when "1000" => HEX <= "0000000"; -- 8
            when "1001" => HEX <= "0010000"; -- 9
            when "1010" => HEX <= "0001000"; -- A
            when "1011" => HEX <= "0000011"; -- B
            when "1100" => HEX <= "1000110"; -- C
            when "1101" => HEX <= "0100001"; -- D
            when "1110" => HEX <= "0000110"; -- E
            when "1111" => HEX <= "0001110"; -- F
            when others => HEX <= "1111111"; -- Apagar display
				
        end case;
    end process;
end Behavioral;
