module Restador(input logic a, b, output logic z);

assign z = a & b;

endmodule 